module rom (input wire [5:0] addr, output reg [7:0] data);
    always @(addr) begin
        case(addr)
            6'b000000: data = 8'b00000000; // mwhahahahaha
            6'b000001: data = 8'b01000101; // E
            6'b000010: data = 8'b01001110; // N
            6'b000011: data = 8'b01000111; // G
            6'b000100: data = 8'b01001001; // I
            6'b000101: data = 8'b01001110; // N
            6'b000110: data = 8'b01000101; // E
            6'b000111: data = 8'b01000101; // E
            6'b001000: data = 8'b01010010; // R
            6'b001001: data = 8'b01001001; // I
            6'b001010: data = 8'b01001110; // N
				6'b001011: data = 8'b01000111; // G
				6'b001100: data = 8'b00100000;
            6'b001101: data = 8'b01000001; // A
            6'b001110: data = 8'b01010011; // S
            6'b001111: data = 8'b01010011; // S
            6'b010000: data = 8'b01001001; // I
            6'b010001: data = 8'b01000111; // G
            6'b010010: data = 8'b01001110; // N
            6'b010011: data = 8'b01001101; // M
            6'b010100: data = 8'b01000101; // E
            6'b010101: data = 8'b01001110; // N
				6'b010110: data = 8'b01010100; // T
				6'b010111: data = 8'b00100000;
            6'b011000: data = 8'b01010011; // S
            6'b011001: data = 8'b01010100; // T
            6'b011010: data = 8'b01010101; // U
            6'b011011: data = 8'b01000100; // D
            6'b011100: data = 8'b01000101; // E
            6'b011101: data = 8'b01001110; // N
				6'b011110: data = 8'b01010100; // T
				6'b011111: data = 8'b00100000;
            6'b100000: data = 8'b01000110; // F
            6'b100001: data = 8'b01010000; // P
            6'b100010: data = 8'b01000111; // G
				6'b100011: data = 8'b01000001; // A
				6'b100100: data = 8'b00100000;
            default: data = 8'b00000000;
        endcase
    end
endmodule
